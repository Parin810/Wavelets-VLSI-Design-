package defs is
constant length : integer:= 2;
constant max_length : integer := 3;
constant sample_length : integer := 2; 
end defs;

